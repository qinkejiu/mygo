module mygo_fifo_i32_d1();
endmodule
module mygo_fifo_i32_d4();
endmodule
module mygo_fifo_i1_d1();
endmodule
