// external fifo
module mygo_fifo_i32_d1();
endmodule
