module main();
endmodule : main
module helper();
endmodule // helper
module mygo_fifo_i32_d1();
endmodule : mygo_fifo_i32_d1
module sentinel();
endmodule // sentinel
